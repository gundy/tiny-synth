function [7:0] synth_note_from_midi_note(
  input [6:0] midi_note;
);
endfunction
